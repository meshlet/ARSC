/// SDRAM controller wrapper
module sdram_control_wrapper (
		input  wire [24:0] address,
		input  wire [1:0]  byteenable_n,
		input  wire        chipselect,
		input  wire [15:0] writedata,
		input  wire        read_n,
		input  wire        write_n,
		output wire [15:0] readdata,
		output wire        readdatavalid,
		output wire        waitrequest,
		input  wire        clk,
		output wire [12:0] dram_addr,
		output wire [1:0]  dram_ba,
		output wire        dram_cas_n,
		output wire        dram_cke,
		output wire        dram_cs_n,
		inout  wire [15:0] dram_dq,
		output wire [1:0]  dram_dqm,
		output wire        dram_ras_n,
		output wire        dram_we_n,
		input  wire        reset_n
	);

	wire    rst_ctrl_reset;
	
	sdram_control sdram_control_unit(
		.clk            (clk),
		.reset_n        (~rst_ctrl_reset),
		.az_addr        (address),
		.az_be_n        (byteenable_n),
		.az_cs          (chipselect),
		.az_data        (writedata),
		.az_rd_n        (read_n),
		.az_wr_n        (write_n),
		.za_data        (readdata),
		.za_valid       (readdatavalid),
		.za_waitrequest (waitrequest),
		.zs_addr        (dram_addr),
		.zs_ba          (dram_ba),
		.zs_cas_n       (dram_cas_n),
		.zs_cke         (dram_cke),
		.zs_cs_n        (dram_cs_n),
		.zs_dq          (dram_dq),
		.zs_dqm         (dram_dqm),
		.zs_ras_n       (dram_ras_n),
		.zs_we_n        (dram_we_n)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),
		.clk            (clk),
		.reset_out      (rst_ctrl_reset),
		.reset_req      (),
		.reset_req_in0  (1'b0),
		.reset_in1      (1'b0),
		.reset_req_in1  (1'b0),
		.reset_in2      (1'b0),
		.reset_req_in2  (1'b0),
		.reset_in3      (1'b0),
		.reset_req_in3  (1'b0),
		.reset_in4      (1'b0),
		.reset_req_in4  (1'b0),
		.reset_in5      (1'b0),
		.reset_req_in5  (1'b0),
		.reset_in6      (1'b0),
		.reset_req_in6  (1'b0),
		.reset_in7      (1'b0),
		.reset_req_in7  (1'b0),
		.reset_in8      (1'b0),
		.reset_req_in8  (1'b0),
		.reset_in9      (1'b0),
		.reset_req_in9  (1'b0),
		.reset_in10     (1'b0),
		.reset_req_in10 (1'b0),
		.reset_in11     (1'b0),
		.reset_req_in11 (1'b0),
		.reset_in12     (1'b0),
		.reset_req_in12 (1'b0),
		.reset_in13     (1'b0),
		.reset_req_in13 (1'b0),
		.reset_in14     (1'b0),
		.reset_req_in14 (1'b0),
		.reset_in15     (1'b0),
		.reset_req_in15 (1'b0)
	);

endmodule
