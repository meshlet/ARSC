//Legal Notice: (C)2017 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

/// ONCHIP MAIN MEMORY
///
/// ARSC system can be configured to use dedicated on-chip memory as its
/// RAM and this chip servers this purpose. It instantiates and configures
/// 64K x 16b of on-chip memory that can be written and read by the ARSC
/// CPU. Additionally, the memory contents can be changed during runtime
/// so that new programs can be loaded without having to re-compile the
/// entire design
module onchip_main_ram
(
	// inputs:
	address,
	byteenable,
	chipselect,
	clk,
	clken,
	reset,
	reset_req,
	write,
	writedata,

	// outputs:
	readdata
);

	parameter INIT_FILE = "arsc_main_memory_init.mif";

	output  [ 15: 0] readdata;
	input   [ 15: 0] address;
	input   [  1: 0] byteenable;
	input            chipselect;
	input            clk;
	input            clken;
	input            reset;
	input            reset_req;
	input            write;
	input   [ 15: 0] writedata;

	wire             clocken0;
	wire    [ 15: 0] readdata;
	wire             wren;
	assign wren = chipselect & write;
	assign clocken0 = clken & ~reset_req;
  
	altsyncram the_altsyncram
    (
		.address_a (address),
		.byteena_a (byteenable),
		.clock0 (clk),
		.clocken0 (clocken0),
		.data_a (writedata),
		.q_a (readdata),
		.wren_a (wren)
	);

	defparam
		the_altsyncram.byte_size = 8,
		the_altsyncram.init_file = INIT_FILE,
		the_altsyncram.lpm_hint = "ENABLE_RUNTIME_MOD=YES, INSTANCE_NAME=ARSC",
		the_altsyncram.lpm_type = "altsyncram",
		the_altsyncram.maximum_depth = 65536,
		the_altsyncram.numwords_a = 65536,
		the_altsyncram.operation_mode = "SINGLE_PORT",
		the_altsyncram.outdata_reg_a = "UNREGISTERED",
		the_altsyncram.ram_block_type = "AUTO",
		the_altsyncram.read_during_write_mode_mixed_ports = "DONT_CARE",
		the_altsyncram.width_a = 16,
		the_altsyncram.width_byteena_a = 2,
		the_altsyncram.widthad_a = 16;

endmodule
